library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Prueba is
    --generic();
    port(
        A : in std_logic_vector(2 downto 0);
        B : out std_logic_vector(2 downto 0);
        );
end entity;

architecture RTL of Prueba is
    
begin
    
end RTL;